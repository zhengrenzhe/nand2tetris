module ThreeWayChoicer(
  a, 
  b, 
  c, 
  out
);
  output out;
  input a;
  input b;
  input c;

endmodule // ThreeWayChoicer